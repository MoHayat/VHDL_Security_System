library ieee;
use ieee.std_logic_1164.all;

entity RAM_tb is
end RAM_tb;

architecture test of RAM_tb is
  -- constants
  constant clk_period : time := 40 ns;

  -- signals
  signal clk_s : std_logic;
  signal n_reset_s      : std_logic;
  signal rd_en_s        : std_logic_vector(2 downto 0);
  signal wr_en_s        : std_logic_vector(2 downto 0);
  signal data_in_s      : std_logic_vector(7 downto 0);
  signal data_out_r_s   : std_logic_vector(7 downto 0);
  signal data_out_g_s   : std_logic_vector(7 downto 0);
  signal data_out_b_s   : std_logic_vector(7 downto 0);
  signal row_s          : integer;
  signal column_s       : integer;

begin

  --instantiate RAM module to begin testing
  RAM_uut : entity work.RAM(hybrid)
  port map(
    clk => clk_s,
    n_reset    => n_reset_s,
    wr_en      => wr_en_s,
    data_in    => data_in_s,
    data_out_r => data_out_r_s,
    data_out_g => data_out_g_s,
    data_out_b => data_out_b_s,
    row        => row_s,
    column     => column_s
  );

  clk_process : process
  begin
    clk_s <= '0';
    wait for clk_period/2;
    clk_s <= '1';
    wait for clk_period/2;
  end process;

  -- stimulus Process
  stim_process : process
  begin
   n_reset_s <= '0';

   wr_en_s   <= "000";

   n_reset_s <= '1';
   wr_en_s   <= "100";
    wait for 40 ns;
   data_in_s <= "00111000";
   wait for 40 ns;
   data_in_s <= "10101011";
   wait for 40 ns;
   data_in_s <= "11110000";
   wait for 40 ns;

   wr_en_s   <= "000";
   wait for 50 ns;

   wr_en_s   <= "010";
   data_in_s <= "00111000";
   wait for 40 ns;
   data_in_s <= "10101011";
   wait for 40 ns;
   data_in_s <= "11110000";
   wait for 40 ns;
   wr_en_s   <= "000";
   wait for 50 ns;

   wr_en_s   <= "001";
   data_in_s <= "00111000";
   wait for 40 ns;
   data_in_s <= "10101011";
   wait for 40 ns;
   data_in_s <= "11110000";
   wait for 40 ns;
   wr_en_s <= "000";
   wait;
   end process;
end test;